red   <= 0;
            green <= 0;
            blue  <= 0;
        end